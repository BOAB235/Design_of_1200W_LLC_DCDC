* NMOS_MODEL_Test1_V2

V3 N001 0 48
V4 N003 0 PULSE(0 10 0 200n 200n 1u 2u)  ; Added pulse width for completeness

R2 N004 N003 3
XM4 N002 N004 0 IRF150P221_L0
XM1 N001 N002 N002 IRF150P221_L0
L1 N001 N002 1u Rser=0.01 Rpar=1Meg Cpar=100p
.tran 1.6u
.include IRF150P221.lib
.ic i(L1)=0
.end
